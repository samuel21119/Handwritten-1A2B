module Character #(
    parameter [9:0] originX = 10'h0,
    parameter [9:0] originY = 10'h0,
    parameter [9:0] width = 10'd40,
    parameter [9:0] height = 10'd80,
    parameter [4:0] characterWidth = 5'd8,
    parameter [4:0] characterHeight = 5'd16
) (
    input [7:0] code,
    input [9:0] h_cnt,
    input [9:0] v_cnt,
    output pixelEnable
);
    localparam [3:0] unitSize = width / characterWidth;

    reg [0:(characterWidth * characterHeight - 1)] flat;

    wire [9:0] clientX = h_cnt - originX;
    wire [9:0] clientY = v_cnt - originY;

    wire [9:0] characterClientX = clientX / unitSize;
    wire [9:0] characterClientY = clientY / unitSize;

    wire valid = (clientX >= 0 && clientX < width) && (clientY >= 0 && clientY < height);
    wire [9:0] index = characterClientX + characterWidth * characterClientY;

    always @(*) begin
        case (code)
            8'h0: begin
                flat = {
                    8'b00111000,
                    8'b01000100,
                    8'b10000010,
                    8'b10000010,
                    8'b10000010,
                    8'b10000010,
                    8'b10000010,
                    8'b10000010,
                    8'b10000010,
                    8'b10000010,
                    8'b10000010,
                    8'b10000010,
                    8'b10000010,
                    8'b10000010,
                    8'b01000100,
                    8'b00111000
                };
            end
            8'h1: begin
                flat = {
                    8'b00001000,
                    8'b00011000,
                    8'b01101000,
                    8'b00001000,
                    8'b00001000,
                    8'b00001000,
                    8'b00001000,
                    8'b00001000,
                    8'b00001000,
                    8'b00001000,
                    8'b00001000,
                    8'b00001000,
                    8'b00001000,
                    8'b00001000,
                    8'b00001000,
                    8'b00001000
                };
            end
            8'h2: begin
                flat = {
                    8'b00111000,
                    8'b01000100,
                    8'b10000010,
                    8'b10000010,
                    8'b10000010,
                    8'b00000010,
                    8'b00000010,
                    8'b00000010,
                    8'b00000010,
                    8'b00000100,
                    8'b00001000,
                    8'b00010000,
                    8'b00100000,
                    8'b01000000,
                    8'b10000000,
                    8'b11111111
                };
            end
            8'h3: begin
                flat = {
                    8'b00111000,
                    8'b01000100,
                    8'b10000010,
                    8'b10000010,
                    8'b10000010,
                    8'b00000010,
                    8'b00000010,
                    8'b00000010,
                    8'b01111100,
                    8'b00000010,
                    8'b00000010,
                    8'b10000010,
                    8'b10000010,
                    8'b10000010,
                    8'b01000100,
                    8'b00111000
                };
            end
            8'h4: begin
                flat = {
                    8'b00000100,
                    8'b00001100,
                    8'b00010100,
                    8'b00010100,
                    8'b00100100,
                    8'b01000100,
                    8'b01000100,
                    8'b10000100,
                    8'b11111110,
                    8'b00000100,
                    8'b00000100,
                    8'b00000100,
                    8'b00000100,
                    8'b00000100,
                    8'b00000100,
                    8'b00000100
                };
            end
            8'h5: begin
                flat = {
                    8'b11111110,
                    8'b10000000,
                    8'b10000000,
                    8'b10000000,
                    8'b10000000,
                    8'b10111000,
                    8'b11000100,
                    8'b10000010,
                    8'b00000010,
                    8'b00000010,
                    8'b00000010,
                    8'b10000010,
                    8'b10000010,
                    8'b10000010,
                    8'b01000100,
                    8'b00111000
                };
            end
            8'h6: begin
                flat = {
                    8'b00111000,
                    8'b01000100,
                    8'b10000010,
                    8'b10000000,
                    8'b10000000,
                    8'b10000000,
                    8'b10000000,
                    8'b10111000,
                    8'b11000100,
                    8'b10000010,
                    8'b10000010,
                    8'b10000010,
                    8'b10000010,
                    8'b10000010,
                    8'b01000100,
                    8'b00111000
                };
            end
            8'h7: begin
                flat = {
                    8'b11111110,
                    8'b10000010,
                    8'b00000010,
                    8'b00000010,
                    8'b00000010,
                    8'b00000010,
                    8'b00000100,
                    8'b00000100,
                    8'b00000100,
                    8'b00001000,
                    8'b00001000,
                    8'b00010000,
                    8'b00010000,
                    8'b00010000,
                    8'b00010000,
                    8'b00010000
                };
            end
            8'h8: begin
                flat = {
                    8'b00111000,
                    8'b01000100,
                    8'b10000010,
                    8'b10000010,
                    8'b10000010,
                    8'b10000010,
                    8'b10000010,
                    8'b01111100,
                    8'b10000010,
                    8'b10000010,
                    8'b10000010,
                    8'b10000010,
                    8'b10000010,
                    8'b10000010,
                    8'b01000100,
                    8'b00111000
                };
            end
            8'h9: begin
                flat = {
                    8'b00111000,
                    8'b01000100,
                    8'b10000010,
                    8'b10000010,
                    8'b10000010,
                    8'b10000010,
                    8'b10000010,
                    8'b01000110,
                    8'b00111010,
                    8'b00000010,
                    8'b00000010,
                    8'b10000010,
                    8'b10000010,
                    8'b10000010,
                    8'b01000100,
                    8'b00111000
                };
            end
            8'ha: begin
                flat = {
                    8'b00000000,
                    8'b00000000,
                    8'b00000000,
                    8'b00000000,
                    8'b00000000,
                    8'b00000000,
                    8'b00000000,
                    8'b00000000,
                    8'b11111100,
                    8'b00000010,
                    8'b00000010,
                    8'b01111110,
                    8'b10000010,
                    8'b10000010,
                    8'b10000010,
                    8'b01111110
                };
            end
            8'hb: begin
                flat = {
                    8'b10000000,
                    8'b10000000,
                    8'b10000000,
                    8'b10000000,
                    8'b10000000,
                    8'b10000000,
                    8'b10000000,
                    8'b10000000,
                    8'b10111000,
                    8'b11000100,
                    8'b10000010,
                    8'b10000010,
                    8'b10000010,
                    8'b10000010,
                    8'b10000100,
                    8'b01111000
                };
            end
            "C": begin
                flat = {
                    8'b00111000,
                    8'b11000100,
                    8'b10000010,
                    8'b10000010,
                    8'b10000000,
                    8'b10000000,
                    8'b10000000,
                    8'b10000000,
                    8'b10000000,
                    8'b10000000,
                    8'b10000000,
                    8'b10000000,
                    8'b10000010,
                    8'b10000010,
                    8'b01000100,
                    8'b00111000
                };
            end
            "E": begin
                flat = {
                    8'b11111110,
                    8'b10000000,
                    8'b10000000,
                    8'b10000000,
                    8'b10000000,
                    8'b10000000,
                    8'b10000000,
                    8'b11111100,
                    8'b10000000,
                    8'b10000000,
                    8'b10000000,
                    8'b10000000,
                    8'b10000000,
                    8'b10000000,
                    8'b10000000,
                    8'b11111110
                };
            end
            "e": begin
                flat = {
                    8'b00000000,
                    8'b00000000,
                    8'b00000000,
                    8'b00000000,
                    8'b00000000,
                    8'b00000000,
                    8'b00000000,
                    8'b00000000,
                    8'b01111100,
                    8'b10000010,
                    8'b10000010,
                    8'b11111110,
                    8'b10000000,
                    8'b10000000,
                    8'b10000010,
                    8'b01111100
                };
            end
            "l": begin
                flat = {
                    8'b00010000,
                    8'b01110000,
                    8'b00010000,
                    8'b00010000,
                    8'b00010000,
                    8'b00010000,
                    8'b00010000,
                    8'b00010000,
                    8'b00010000,
                    8'b00010000,
                    8'b00010000,
                    8'b00010000,
                    8'b00010000,
                    8'b00010000,
                    8'b00010000,
                    8'b11111110
                };
            end
            "n": begin
                flat = {
                    8'b00000000,
                    8'b00000000,
                    8'b00000000,
                    8'b00000000,
                    8'b00000000,
                    8'b00000000,
                    8'b00000000,
                    8'b00000000,
                    8'b10011000,
                    8'b10100100,
                    8'b11000010,
                    8'b10000010,
                    8'b10000010,
                    8'b10000010,
                    8'b10000010,
                    8'b10000010
                };
            end
            "r": begin
                flat = {
                    8'b00000000,
                    8'b00000000,
                    8'b00000000,
                    8'b00000000,
                    8'b00000000,
                    8'b00000000,
                    8'b00000000,
                    8'b00000000,
                    8'b10011100,
                    8'b10100010,
                    8'b11000000,
                    8'b10000000,
                    8'b10000000,
                    8'b10000000,
                    8'b10000000,
                    8'b10000000
                };
            end
            "t": begin
                flat = {
                    8'b10000000,
                    8'b10000000,
                    8'b10000000,
                    8'b10000000,
                    8'b10000000,
                    8'b11111110,
                    8'b10000000,
                    8'b10000000,
                    8'b10000000,
                    8'b10000000,
                    8'b10000000,
                    8'b10000000,
                    8'b10000000,
                    8'b10000000,
                    8'b01000010,
                    8'b00111100
                };
            end
            default: begin
                flat = {
                    8'b00000000,
                    8'b00000000,
                    8'b00000000,
                    8'b00000000,
                    8'b00000000,
                    8'b00000000,
                    8'b00000000,
                    8'b00000000,
                    8'b00000000,
                    8'b00000000,
                    8'b00000000,
                    8'b00000000,
                    8'b00000000,
                    8'b00000000,
                    8'b00000000,
                    8'b00000000
                };
            end
        endcase
    end

    // only output pixel when showing character
    assign pixelEnable = valid & flat[index];

endmodule